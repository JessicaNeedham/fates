CDF       
      
fates_NCWD        fates_history_age_bins        fates_history_height_bins         fates_history_size_bins    (   fates_hydr_organs         fates_leafage_class       fates_litterclass         	fates_pft         fates_prt_organs      fates_scalar      fates_string_length    <   fates_variants              history       �This file was made from FatesPFTIndexSwapper.py 
 Input File = parameter_files/fates_params_Ssenes_default.nc 
 Indices = [1, 1]      �   !fates_history_sizeclass_bin_edges                  units         cm     	long_name         OLower edges for DBH size class bins used in size-resolved cohort history output       �  w�    fates_history_ageclass_bin_edges               units         yr     	long_name         HLower edges for age class bins used in age-resolved patch history output        xL   fates_prt_organ_name         
         units         unitless - string      	long_name         5Plant organ name (order must match PRTGenericMod.F90)        h  xh   fates_prt_alloc_priority                  units         index (0-fates_prt_organs)     	long_name         Priority order for allocation         0  y�   fates_prt_nitr_stoich_p1                  units         (gN/gC)    	long_name         #nitrogen stoichiometry, parameter 1       0  z    fates_prt_nitr_stoich_p2                  units         (gN/gC)    	long_name         #nitrogen stoichiometry, parameter 2       0  z0   fates_prt_phos_stoich_p1                  units         (gP/gC)    	long_name         &phosphorous stoichiometry, parameter 1        0  z`   fates_prt_phos_stoich_p2                  units         (gP/gC)    	long_name         &phosphorous stoichiometry, parameter 2        0  z�   fates_turnover_carb_retrans                   units         -      	long_name         .retranslocation fraction of carbon in turnover        0  z�   fates_turnover_nitr_retrans                   units         -      	long_name         0retranslocation fraction of nitrogen in turnover      0  z�   fates_turnover_phos_retrans                   units         -      	long_name         @retranslocation fraction of phosphorous in turnover, parameter 1      0  {    	fates_FBD                  units         NA     	long_name         ?spitfire parameter related to fuel bulk density, see SFMain.F90         {P   	fates_SAV                  units         NA     	long_name         Jspitfire parameter related to surface area to volume ratio, see SFMain.F90          {h   fates_history_height_bin_edges                 units         m      	long_name         BLower edges for height bins used in height-resolved history output          {�   fates_low_moisture_Coeff               units         NA     	long_name         3spitfire parameter, equation B1 Thonicke et al 2010         {�   fates_low_moisture_Slope               units         NA     	long_name         3spitfire parameter, equation B1 Thonicke et al 2010         {�   fates_max_decomp               units         kgC/m2/yr ?    	long_name         Wmaximum rate of litter & CWD transfer from non-decomposing class into decomposing class         {�   fates_mid_moisture                 units         NA     	long_name         >spitfire litter moisture threshold to be considered medium dry          {�   fates_mid_moisture_Coeff               units         NA     	long_name         3spitfire parameter, equation B1 Thonicke et al 2010         {�   fates_mid_moisture_Slope               units         NA     	long_name         3spitfire parameter, equation B1 Thonicke et al 2010         |   fates_min_moisture                 units         NA     	long_name         <spitfire litter moisture threshold to be considered very dry        |(   fates_hydr_avuln_node                     units         unitless   	long_name         )xylem vulnerability curve shape parameter            |@   fates_hydr_epsil_node                     units         MPa    	long_name         bulk elastic modulus         |`   fates_hydr_fcap_node                  units         unitless   	long_name         6fraction of (1-resid_node) that is capillary in source           |�   fates_hydr_kmax_node                  units         	kgMPa/m/s      	long_name         9maximum xylem conductivity per unit conducting xylem area            |�   fates_hydr_p50_node                   units         MPa    	long_name         1xylem water potential at 50% loss of conductivity            |�   fates_hydr_pinot_node                     units         MPa    	long_name          osmotic potential at full turgor         |�   fates_hydr_pitlp_node                     units         MPa    	long_name         turgor loss point            }    fates_hydr_resid_node                     units         fraction   	long_name         residual fraction            }    fates_hydr_thetas_node                    units         cm3/cm3    	long_name         saturated water content          }@   fates_CWD_frac                  units         fraction   	long_name         ;fraction of woody (bdead+bsw) biomass destined for CWD pool         }`   fates_pftname            
         units         unitless - string      	long_name         Description of plant type         x  }p   fates_rootprof_beta                   units         unitless   	long_name         QRooting beta parameter, for C and N vertical discretization (NOT USED BY DEFAULT)           }�   fates_alloc_storage_cushion                units         fraction   	long_name         Gmaximum size of storage C pool, relative to maximum size of leaf C pool         }�   fates_allom_agb1               units         variable   	long_name         Parameter 1 for agb allometry           ~    fates_allom_agb2               units         variable   	long_name         Parameter 2 for agb allometry           ~   fates_allom_agb3               units         variable   	long_name         Parameter 3 for agb allometry           ~   fates_allom_agb4               units         variable   	long_name         Parameter 4 for agb allometry           ~   fates_allom_agb_frac               units         fraction   	long_name         .Fraction of woody biomass that is above ground          ~    fates_allom_amode                  units         index      	long_name         AGB allometry function index        ~(   fates_allom_blca_expnt_diff                units         unitless   	long_name         Ddifference between allometric DBH:bleaf and DBH:crown area exponents        ~0   fates_allom_cmode                  units         index      	long_name         ,coarse root biomass allometry function index        ~8   fates_allom_d2bl1                  units         variable   	long_name         Parameter 1 for d2bl allometry          ~@   fates_allom_d2bl2                  units         variable   	long_name         Parameter 2 for d2bl allometry          ~H   fates_allom_d2bl3                  units         unitless   	long_name         Parameter 3 for d2bl allometry          ~P    fates_allom_d2ca_coefficient_max               units         m2 cm^(-1/beta)    	long_name         Omax (savanna) dbh to area multiplier factor where: area = n*d2ca_coeff*dbh^beta         ~X    fates_allom_d2ca_coefficient_min               units         m2 cm^(-1/beta)    	long_name         Nmin (forest) dbh to area multiplier factor where: area = n*d2ca_coeff*dbh^beta          ~`   fates_allom_d2h1               units         variable   	long_name         /Parameter 1 for d2h allometry (intercept, or c)         ~h   fates_allom_d2h2               units         variable   	long_name         +Parameter 2 for d2h allometry (slope, or m)         ~p   fates_allom_d2h3               units         variable   	long_name         (Parameter 3 for d2h allometry (optional)        ~x   fates_allom_dbh_maxheight                  units         cm     	long_name         Ythe diameter (if any) corresponding to maximum height, diameters may increase beyond this           ~�   fates_allom_fmode                  units         index      	long_name         *fine root biomass allometry function index          ~�   fates_allom_frbstor_repro                  units         fraction   	long_name         8fraction of bstore goes to reproduction after plant dies        ~�   fates_allom_hmode                  units         index      	long_name         height allometry function index         ~�   fates_allom_l2fr               units         gC/gC      	long_name         ,Allocation parameter: fine root C per leaf C        ~�   fates_allom_la_per_sa_int                  units         m2/cm2     	long_name         %Leaf area per sapwood area, intercept           ~�   fates_allom_la_per_sa_slp                  units         m2/cm2/m   	long_name         GLeaf area per sapwood area rate of change with height, slope (optional)         ~�   fates_allom_lmode                  units         index      	long_name         %leaf biomass allometry function index           ~�   fates_allom_sai_scaler                 units         m2/m2      	long_name         allometric ratio of SAI per LAI         ~�   fates_allom_smode                  units         index      	long_name          sapwood allometry function index        ~�   fates_allom_stmode                 units         index      	long_name          storage allometry function index        ~�   fates_branch_turnover                  units         yr-1   	long_name         turnover time of branches           ~�   	fates_c2b                  units         ratio      	long_name         7Carbon to biomass multiplier of bulk structural tissues         ~�   fates_displar                  units         unitless   	long_name         1Ratio of displacement height to canopy top height           ~�   fates_fire_alpha_SH                units         NA     	long_name         Hspitfire parameter, alpha scorch height, Equation 16 Thonicke et al 2010        ~�   fates_fire_bark_scaler                 units         fraction   	long_name         8the thickness of a cohorts bark as a fraction of its dbh        ~�   fates_fire_crown_depth_frac                units         fraction   	long_name         8the depth of a cohorts crown as a fraction of its height            fates_fire_crown_kill                  units         NA     	long_name         6fire parameter, see equation 22 in Thonicke et al 2010             fates_fr_fcel                  units         fraction   	long_name         #Fine root litter cellulose fraction            fates_fr_flab                  units         fraction   	long_name          Fine root litter labile fraction           fates_fr_flig                  units         fraction   	long_name          Fine root litter lignin fraction            fates_grperc               units         unitless   	long_name         Growth respiration factor           (   fates_hydr_avuln_gs                units         unitless   	long_name         @shape parameter for stomatal control of water vapor exiting leaf        0   fates_hydr_p50_gs                  units         MPa    	long_name         3water potential at 50% loss of stomatal conductance         8   fates_hydr_p_taper                 units         unitless   	long_name         xylem taper exponent        @   fates_hydr_rfrac_stem                  units         fraction   	long_name         6fraction of total tree resistance from troot to canopy          H   fates_hydr_rs2                 units         m      	long_name         absorbing root radius           P   fates_hydr_srl                 units         m g-1      	long_name         specific root length        X   fates_leaf_BB_slope                units         unitless   	long_name         +stomatal slope parameter, as per Ball-Berry         `   fates_leaf_c3psn               units         flag   	long_name         #Photosynthetic pathway (1=c3, 0=c4)         h   fates_leaf_clumping_index                  units         fraction (0-1)     	long_name         bfactor describing how much self-occlusion of leaf scattering elements decreases light interception          p   fates_leaf_diameter                units         m      	long_name         Characteristic leaf dimension           x   fates_leaf_jmaxha                  units         J/mol      	long_name         activation energy for jmax          �   fates_leaf_jmaxhd                  units         J/mol      	long_name         deactivation energy for jmax        �   fates_leaf_jmaxse                  units         J/mol/K    	long_name         entropy term for jmax           �   fates_leaf_slamax                  units         m^2/gC     	long_name         >Maximum Specific Leaf Area (SLA), even if under a dense canopy          �   fates_leaf_slatop                  units         m^2/gC     	long_name         ?Specific Leaf Area (SLA) at top of canopy, projected area basis         �   fates_leaf_stor_priority               units         unitless   	long_name         7factor governing priority of replacing storage with NPP         �   fates_leaf_tpuha               units         J/mol      	long_name         activation energy for tpu           �   fates_leaf_tpuhd               units         J/mol      	long_name         deactivation energy for tpu         �   fates_leaf_tpuse               units         J/mol/K    	long_name         entropy term for tpu        �   fates_leaf_vcmaxha                 units         J/mol      	long_name         activation energy for vcmax         �   fates_leaf_vcmaxhd                 units         J/mol      	long_name         deactivation energy for vcmax           �   fates_leaf_vcmaxse                 units         J/mol/K    	long_name         entropy term for vcmax          �   fates_leaf_xl                  units         unitless   	long_name         Leaf/stem orientation index         �   fates_lf_fcel                  units         fraction   	long_name         Leaf litter cellulose fraction          �   fates_lf_flab                  units         fraction   	long_name         Leaf litter labile fraction         �   fates_lf_flig                  units         fraction   	long_name         Leaf litter lignin fraction         �   #fates_maintresp_reduction_curvature                units         unitless (0-1)     	long_name         Gcurvature of MR reduction as f(carbon storage), 1=linear, 0=very curved         �    #fates_maintresp_reduction_intercept                units         unitless (0-1)     	long_name         Qintercept of MR reduction as f(carbon storage), 0=no throttling, 1=max throttling           �   fates_mort_bmort               units         1/yr   	long_name         background mortality rate           �   fates_mort_freezetol               units         NA     	long_name         (minimum temperature tolerance (NOT USED)        �   fates_mort_hf_flc_threshold                units         fraction   	long_name         [plant fractional loss of conductivity at which drought mortality begins for hydraulic model         �    fates_mort_hf_sm_threshold                 units         unitless   	long_name         Usoil moisture (btran units) at which drought mortality begins for non-hydraulic model           �(   fates_mort_ip_senescence               units         dbh cm     	long_name         %Mortality senescence inflection point           �0   fates_mort_r_senescence                units         mortality rate dbh^-1      	long_name         #Mortality senescence rate of change         �8   fates_mort_scalar_coldstress               units         1/yr   	long_name         'maximum mortality rate from cold stress         �@   fates_mort_scalar_cstarvation                  units         1/yr   	long_name         -maximum mortality rate from carbon starvation           �H   fates_mort_scalar_hydrfailure                  units         1/yr   	long_name         -maximum mortality rate from hydraulic failure           �P   fates_pft_used                 units          0 = off (dont use), 1 = on (use)   	long_name         DSwitch to turn on and off PFTs (also see fates_initd for cold-start)        �X   fates_phen_evergreen               units         logical flag   	long_name         $Binary flag for evergreen leaf habit        �`   fates_phen_season_decid                units         logical flag   	long_name         -Binary flag for seasonal-deciduous leaf habit           �h   fates_phen_stress_decid                units         logical flag   	long_name         +Binary flag for stress-deciduous leaf habit         �p   fates_phenflush_fraction               units         fraction   	long_name         OUpon bud-burst, the maximum fraction of storage carbon used for flushing leaves         �x   !fates_prescribed_mortality_canopy                  units         1/yr   	long_name         =mortality rate of canopy trees for prescribed physiology mode           ��   %fates_prescribed_mortality_understory                  units         1/yr   	long_name         Amortality rate of understory trees for prescribed physiology mode           ��   fates_prescribed_npp_canopy                units         gC / m^2 / yr      	long_name         FNPP per unit crown area of canopy trees for prescribed physiology mode          ��   fates_prescribed_npp_understory                units         gC / m^2 / yr      	long_name         JNPP per unit crown area of understory trees for prescribed physiology mode          ��   fates_prescribed_recruitment               units         n/yr   	long_name         /recruitment rate for prescribed physiology mode         ��   fates_recruit_hgt_min                  units         m      	long_name         Bthe minimum height (ie starting height) of a newly recruited plant          ��   fates_recruit_initd                units         stems/m2   	long_name         Einitial seedling density for a cold-start near-bare-ground simulation           ��   fates_rholnir                  units         fraction   	long_name         Leaf reflectance: near-IR           ��   fates_rholvis                  units         fraction   	long_name         Leaf reflectance: visible           ��   fates_rhosnir                  units         fraction   	long_name         Stem reflectance: near-IR           ��   fates_rhosvis                  units         fraction   	long_name         Stem reflectance: visible           ��   fates_root_long                units         yr     	long_name         -root longevity (alternatively, turnover time)           ��   fates_roota_par                units         1/m    	long_name         "CLM rooting distribution parameter          ��   fates_rootb_par                units         1/m    	long_name         "CLM rooting distribution parameter          ��   fates_seed_alloc               units         fraction   	long_name         7fraction of available carbon balance allocated to seeds         ��   fates_seed_alloc_mature                units         fraction   	long_name         cfraction of available carbon balance allocated to seeds in mature plants (adds to fates_seed_alloc)         ��   fates_seed_dbh_repro_threshold                 units         cm     	long_name         Ythe diameter (if any) where the plant will start extra clonal allocation to the seed pool           �    fates_seed_decay_turnover                  units         1/yr   	long_name         3turnover time for seeds with respect to germination         �    fates_seed_germination_timescale               units         1/yr   	long_name         -turnover time for seeds with respect to decay           �   fates_seed_rain                units         	KgC/m2/yr      	long_name         :External seed rain from outside site (non-mass conserving)          �   fates_senleaf_long_fdrought                units         unitless[0-1]      	long_name         Kmultiplication factor for leaf longevity of senescent leaves during drought         �    fates_smpsc                units         mm     	long_name         -Soil water potential at full stomatal closure           �(   fates_smpso                units         mm     	long_name         -Soil water potential at full stomatal opening           �0   fates_taulnir                  units         fraction   	long_name         Leaf transmittance: near-IR         �8   fates_taulvis                  units         fraction   	long_name         Leaf transmittance: visible         �@   fates_tausnir                  units         fraction   	long_name         Stem transmittance: near-IR         �H   fates_tausvis                  units         fraction   	long_name         Stem transmittance: visible         �P   fates_trim_inc                 units         m2/m2      	long_name         2Arbitrary incremental change in trimming function.          �X   fates_trim_limit               units         m2/m2      	long_name         6Arbitrary limit to reductions in leaf area with stress          �`   fates_turnover_retrans_mode                units         index      	long_name         1retranslocation method for leaf/fineroot turnover           �h   fates_wood_density                 units         g/cm3      	long_name         %mean density of woody tissue in plant           �p   fates_woody                units         logical flag   	long_name         Binary woody lifeform flag          �x   
fates_z0mr                 units         unitless   	long_name         7Ratio of momentum roughness length to canopy top height         ��   fates_leaf_long                   units         yr     	long_name         &Leaf longevity (ie turnover timescale)          ��   fates_leaf_vcmax25top                     units         umol CO2/m^2/s     	long_name         5maximum carboxylation rate of Rub. at 25C, canopy top           ��   fates_base_mr_20      	         units         gC/gN/s    	long_name         DBase maintenance respiration rate for plant tissues, using Ryan 1991        ��   fates_bbopt_c3        	         units         umol H2O/m**2/s    	long_name         5Ball-Berry minimum unstressed leaf conductance for C3           ��   fates_bbopt_c4        	         units         umol H2O/m**2/s    	long_name         5Ball-Berry minimum unstressed leaf conductance for C4           ��   fates_canopy_closure_thresh       	         units         unitless   	long_name         Wtree canopy coverage at which crown area allometry changes from savanna to forest value         ��   fates_cohort_fusion_tol       	         units         unitless   	long_name         5minimum fraction in difference in dbh between cohorts           ��   fates_comp_excln      	         units         none   	long_name         Kweighting factor (exponent on dbh) for canopy layer exclusion and promotion         ��   fates_cwd_fcel        	         units         unitless   	long_name         Cellulose fraction for CWD          ��   fates_cwd_flig        	         units         unitless   	long_name         &Lignin fraction of coarse woody debris          ��   fates_fire_nignitions         	         units         /m2 (?)    	long_name         @number of daily ignitions (nfires = nignitions*FDI*area_scaling)        ��   fates_hydr_kmax_rsurf         	         units         kg water/m2 root area/Mpa/s    	long_name         +maximum conducitivity for unit root surface         ��   fates_hydr_psi0       	         units         MPa    	long_name         %sapwood water potential at saturation           ��   fates_hydr_psicap         	         units         MPa    	long_name         =sapwood water potential at which capillary reserves exhausted           ��   fates_init_litter         	         units         NA     	long_name         =Initialization value for litter pool in cold-start (NOT USED)           ��   fates_logging_coll_under_frac         	         units         fraction   	long_name         MFraction of stems killed in the understory when logging generates disturbance           ��   fates_logging_collateral_frac         	         units         fraction   	long_name         MFraction of large stems in upperstory that die from logging collateral damage           ��   fates_logging_dbhmax_infra        	         units         cm     	long_name         [Tree diameter, above which infrastructure from logging does not impact damage or mortality.         ��   fates_logging_dbhmin      	         units         cm     	long_name         'Minimum dbh at which logging is applied         ��   fates_logging_direct_frac         	         units         fraction   	long_name         +Fraction of stems logged directly per event         ��   fates_logging_event_code      	         units         unitless   	long_name         ;Integer code that options how logging events are structured         ��   fates_logging_mechanical_frac         	         units         fraction   	long_name         EFraction of stems killed due infrastructure an other mechanical means           ��   fates_mort_disturb_frac       	         units         fraction   	long_name         ffraction of canopy mortality that results in disturbance (i.e. transfer of area from new to old patch)          ��   fates_mort_understorey_death      	         units         fraction   	long_name         Ifraction of plants in understorey cohort impacted by overstorey tree-fall           ��   fates_patch_fusion_tol        	         units         unitless   	long_name         :minimum fraction in difference in profiles between patches          ��   fates_phen_a      	         units         none   	long_name         LGDD accumulation function, intercept parameter: gdd_thesh = a + b exp(c*ncd)        ��   fates_phen_b      	         units         none   	long_name         MGDD accumulation function, multiplier parameter: gdd_thesh = a + b exp(c*ncd)           ��   fates_phen_c      	         units         none   	long_name         KGDD accumulation function, exponent parameter: gdd_thesh = a + b exp(c*ncd)         ��   fates_phen_chiltemp       	         units         	degrees C      	long_name         chilling day counting threshold         �    fates_phen_coldtemp       	         units         	degrees C      	long_name         Ctemperature exceedance to flag a cold-day for temperature leaf drop         �   fates_phen_doff_time      	         units         days   	long_name         Eday threshold compared against days since leaves became off-allometry           �   fates_phen_drought_threshold      	         units         m3/m3      	long_name         =liquid volume in soil layer, threashold for drought phenology           �   fates_phen_mindayson      	         units         days   	long_name         Dday threshold compared against days since leaves became on-allometry        �   fates_phen_ncolddayslim       	         units         days   	long_name         2day threshold exceedance for temperature leaf-drop          �   fates_soil_salinity       	         units         ppt    	long_name         Fsoil salinity used for model when not coupled to dynamic soil salinity          �   fates_drying_ratio               units         NA     	long_name         [spitfire parameter, fire drying ratio for fuel moisture, alpha_FMC EQ 6 Thonicke et al 2010         �   fates_durat_slope                units         NA     	long_name         Lspitfire parameter, fire max duration slope, Equation 14 Thonicke et al 2010        �    fates_fdi_a              units         NA     	long_name         spitfire parameter (unknown)            �$   fates_fdi_alpha              units         NA     	long_name         Wspitfire parameter, EQ 7 Venevsky et al. GCB 2002,(modified EQ 8 Thonicke et al. 2010)          �(   fates_fdi_b              units         NA     	long_name         spitfire parameter (unknown)            �,   fates_fuel_energy                units         kJ/kg      	long_name         'pitfire parameter, heat content of fuel         �0   fates_max_durat              units         minutes    	long_name         Jspitfire parameter, fire maximum duration, Equation 14 Thonicke et al 2010          �4   fates_miner_damp             units         NA     	long_name         Lspitfire parameter, mineral-dampening coefficient EQ A1 Thonicke et al 2010         �8   fates_miner_total                units         fraction   	long_name         Gspitfire parameter, total mineral content, Table A1 Thonicke et al 2010         �<   fates_part_dens              units         kg/m2      	long_name         Kspitfire parameter, oven dry particle density, Table A1 Thonicke et al 2010         �@    @�  A   Ap  A�  A�  A�  B  B   B4  BH  B\  Bp  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  C  C  C  C  C  C  C   C%  C*  C/  C4  C9  C>  CH      ?�  @   @�  A   A�  BH  leaf                                                        fine root                                                   sapwood                                                     storage                                                     reproduction                                                structure                                                   |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  =+=+<ě�<ě�2+�w2+�w2+�w2+�w        ;�u;�u|�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  <���<���                                        |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  |�  AvffA�ffA���Dy� @�  @�  AP  @e�?z�H>L��B�  B�      =���>���?�  @@  A   ?�\)?��?z�H?L��?�33?�33?�R?8Q�?Y��?L��?�R?�R?�>��>��>B�\?�  Dy� ?8Q�?�\>\?�  ?L��?L��@ff?�(�?��?L��@L��@L��@ff?�(�?��?L��@L��@L��>8Q�=�        >u>u@   @   @   @   @   @   @   @   A@  A@  A   A   A   A   A   A           =��
=��
=��
=��
        �y� �y� @@  @@  �y� �y� �y� �y� �  �  �  �  �  �  �  �  ���]���]��1f��1f��1f��1f��������������33��33��33��33��������>�  >�  >�ff>�ff>�ff>�ff>��>��?&ff?&ff?&ff?&ff?&ff?&ff?@  ?@  =8Q�=���>W
=?+�broadleaf_evergreen_tropical_tree                           broadleaf_evergreen_tropical_tree                           ?y�#?y�#|�  |�  ?���?���=�:�=�:�?n�?n�?�Q�?�Q�?nV?nV?��?��?�  ?�          ?�  ?�  =�\)=�\)?�ff?�ff?��?��?('?('>�>�?#�
?#�
>�p�>�p��y���y��B�  B�  ?�  ?�          ?�  ?�  ?�  ?�  ?L��?L��        ?�  ?�  =���=���?�  ?�  ?�  ?�  C  C  @   @   ?+�?+�>L��>L��=�\)=�\)?   ?   ?Fff?Fff?   ?   >�  >�  >�  >�  =�G�=�G�@   @   ��  ��  >�~�>�~�?   ?   8ѷ8ѷA�  A�  A   A   ?�  ?�  ?Y��?Y��=#�
=#�
G* G* Hz Hz C�� C�� =�a=�a<D��<D��?L��?L��GOl GOl H�H�C�  C�  G2 G2 H��H��C� C� =���=���?   ?   >�  >�  >�  >�  <#�
<#�
?�  ?�  <e`B<e`B@   @   ?   ?   5�7�5�7�B�  B�  >L��>L��@@  @@  ?��?��?��?��?�  ?�  ?�  ?�                  |�  |�  <���<���<���<���>���>���=   =   <��
<��
?�ff?�ff>L��>L��>�ff>�ff=���=���>Ǯ>Ǯ>#�
>#�
?�  ?�  @�  @�  ?�  ?�  =���=���        C  C  ?�\?�\?   ?           ?�  ?�  �y �y ǀ� ǀ� >�  >�  =L��=L��:�o:�o:�o:�o<�<�>���>���?�  ?�  ?333?333?�  ?�  =aG�=aG�?�  ?�  BH  BH  6)EF@ G@ ?L��=��
@@  ?B�\>uAp  A�      ���=L��?Q=L��B  BH  >����  =L��?�  ?Q=L��  D� �#�
@�  @�  B�  >��A�  @�  >���FK  �0��A���9���Cs�F�� Cp  >մ$=aG�D @ 